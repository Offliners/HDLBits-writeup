module top_module (
    input clk,
    input reset,      // Synchronous reset
    input data,
    output shift_ena,
    output counting,
    input done_counting,
    output done,
    input ack );
    
    parameter [2:0] IDLE = 3'd0, S0	= 3'd1, S1 = 3'd2, S2 = 3'd3, S3 = 3'd4, SHIFT = 3'd5, COUNT = 3'd6, DONE = 3'd7; 
    reg [3:0] state, next_state;
    reg [2:0] count;
    
    always @(posedge clk) begin
        if (reset) begin
            state <= IDLE;
            count <= 3'd0;
        end
		else begin
            if(state == SHIFT)
                count <= count + 3'd1;
            else
                count <= 3'd1;
                
            state <= next_state;
        end
	end

	always @(*) begin
		case (state) 
            IDLE : next_state <= data ? S1 : IDLE;
            S1 : next_state <= data ? S2 : IDLE;
            S2 : next_state <= data ? S2 : S3;
			S3  : next_state <= data ? SHIFT : IDLE;
            SHIFT : next_state <= count == 3'd4 ? COUNT : SHIFT;
			COUNT : next_state <= done_counting ? DONE : COUNT;
			DONE  : next_state <= ack ? IDLE : DONE;			
		endcase
	end

	assign shift_ena = state == SHIFT;
	assign counting = state == COUNT;
	assign done = state == DONE;

endmodule