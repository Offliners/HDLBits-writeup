module top_module(
    input clk,
    input reset,    // Synchronous reset
    input in,
    output disc,
    output flag,
    output err);
    
    parameter IDLE=0, RECEIVE=1, DISCARD=2, FLAG=3, ERROR=4;
    reg [2:0] state, next_state;
    reg [31:0] count;
    
    always @(posedge clk) begin
        if(reset) begin
            state <= IDLE;
            count <= 0;
        end
        else begin
            if(in)
                count <= count + 1;
            else
                count <= 0;
            
            state <= next_state;
        end
    end
    
    always @(*) begin
        case(state)
            IDLE : next_state <= in ? RECEIVE : IDLE;
            RECEIVE : begin
                case(count)
                    3'd5 : next_state <= in ? RECEIVE : DISCARD;
                    3'd6 : next_state <= in ? ERROR : FLAG;
                    default: next_state <= in ? RECEIVE : IDLE;
                endcase
            end
            DISCARD : next_state <= in ? RECEIVE : IDLE;
            FLAG : next_state <= in ? RECEIVE : IDLE;
            ERROR : next_state <= in ? ERROR : IDLE;
        endcase
    end
    
    assign disc = state == DISCARD;
    assign flag = state == FLAG;
    assign err = state == ERROR;

endmodule
