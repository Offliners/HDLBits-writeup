module top_module (
    input clk,
    input reset,      // Synchronous reset
    input data,
    output reg [3:0] count,
    output counting,
    output done,
    input ack );
    
        parameter [2:0] IDLE = 3'd0, S0	= 3'd1, S1 = 3'd2, S2 = 3'd3, S3 = 3'd4, SHIFT = 3'd5, COUNT = 3'd6, DONE = 3'd7; 
    reg [3:0] state, next_state;
    reg [2:0] shitf_count;
    reg [9:0] count_1k;
    
    always @(posedge clk) begin
        if (reset) begin
            state <= IDLE;
            shitf_count <= 3'd0;
        end
		else begin
            if(state == SHIFT)
                shitf_count <= shitf_count + 3'd1;
            else
                shitf_count <= 3'd1;
                
            state <= next_state;
        end
	end
    
    always @(posedge clk) begin
		case (state) 
            SHIFT : count[3'd4 - shitf_count] <= data;
			COUNT : begin
				if (count >= 0) begin
                    if (count_1k < 10'd999) 
						count_1k <= count_1k + 10'd1;
					else begin
						count <= count - 4'b1;
						count_1k <= 10'd0;
					end
				end
			end
			default : count_1k <= 10'd0;
		endcase
	end

	always @(*) begin
		case (state) 
            IDLE : next_state <= data ? S1 : IDLE;
            S1 : next_state <= data ? S2 : IDLE;
            S2 : next_state <= data ? S2 : S3;
			S3  : next_state <= data ? SHIFT : IDLE;
            SHIFT : next_state <= shitf_count == 3'd4 ? COUNT : SHIFT;
            COUNT : next_state <= (count == 0 && count_1k == 10'd999) ? DONE : COUNT;
			DONE  : next_state <= ack ? IDLE : DONE;			
		endcase
	end

	assign counting = state == COUNT;
	assign done = state == DONE;

endmodule
