module top_module(
    input clk,
    input in,
    input reset,    // Synchronous reset
    output done
); 
    parameter IDLE=0, START=1, STOP=2, ERROR=3;
    reg [1:0] state, next_state;
    reg [3:0] count;
    
    always @(posedge clk) begin
        if(reset) begin
            state <= IDLE;
            count <= 4'b0;
        end
        else begin
            if(state == START && count != 8)
                count <= count + 4'b1;
            else if(state == STOP || state == ERROR)
                count <= 4'b0;
            else
                count <= count;
            
            state <= next_state;
        end
    end
    
    always @(*) begin
        case(state)
            IDLE : next_state <= in ? IDLE : START;
            START : next_state <= (count == 8) ? (in ? STOP : ERROR) : START;
            STOP : next_state <= in ? IDLE : START;
            ERROR : next_state <= in ? IDLE : ERROR;
            default: next_state <= IDLE;
        endcase
    end
    
    assign done = state == STOP;

endmodule