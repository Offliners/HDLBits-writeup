module top_module(
    input clk,
    input in,
    input reset,    // Synchronous reset
    output [7:0] out_byte,
    output done
); //
    parameter IDLE=0, START=1, STOP=2, ERROR=3;
    reg [1:0] state, next_state;
    reg [3:0] count;
    reg [7:0] data;

    // Use FSM from Fsm_serial
    always @(posedge clk) begin
        if(reset) begin
            state <= IDLE;
            count <= 4'b0;
        end
        else begin
            if(state == START && count != 8) begin
                count <= count + 4'b1;
                data <= {in, data[7:1]};
            end
            else if(state == STOP || state == ERROR)
                count <= 4'b0;
            else
                count <= count;
            
            state <= next_state;
        end
    end
    
    always @(*) begin
        case(state)
            IDLE : next_state <= in ? IDLE : START;
            START : next_state <= count == 8 ? (in ? STOP : ERROR) : START;
            STOP : next_state <= in ? IDLE : START;
            ERROR : next_state <= in ? IDLE : ERROR; 
        endcase
    end

    // New: Datapath to latch input bits.
    assign done = state == STOP;
    assign out_byte = done ? data : 8'b0;

endmodule